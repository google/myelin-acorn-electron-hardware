
module internal_osc (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
