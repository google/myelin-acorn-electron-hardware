module bus_scope_main(
	output wire [31:0] fx3_D
);

assign fx3_D = 32'bZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;

endmodule
