-- Copyright 2017 Google Inc.
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cpu_socket_expansion is
    Port (
      -- Buffer chips:

      -- *buf_ext_to_cpu buffers from pins A->B when 1, B->A when 0.
      -- A = pins 2-9, B = pins 18-11.
      -- A pins all connect to the external connector, and B pins connect to
      -- the CPU socket, so setting *buf_ext_to_cpu=0 means the CPU drives the
      -- external port, and setting it to 1 means the external port is driving,
      -- and defaulting to 0 is the most sensible.

      -- *buf_nCE enables buffers when 0, disables when 1.  Defaulting to just
      -- disabling all buffers.

      abuf_ext_to_cpu : out std_logic := '0';
      abuf_nCE : out std_logic := '1';

      dbuf_ext_to_cpu : out std_logic := '0';
      dbuf_nCE : out std_logic := '1';

      -- For shadow RAM support, we buffer A13:A15.  When shadow RAM is not being accessed,
      -- these should just pass through from the CPU to the motherboard.
      cpu_A13_1 : out std_logic; -- connects to motherboard
      cpu_A13_2 : in std_logic; -- connects to ABUFH and socketed CPU
      cpu_A14_1 : out std_logic; -- connects to motherboard
      cpu_A14_2 : in std_logic; -- connects to ABUFH and socketed CPU
      cpu_A15_1 : out std_logic; -- connects to motherboard
      cpu_A15_2 : in std_logic; -- connects to ABUFH and socketed CPU

      -- This may or may not connect to the ULA's 16MHz clock; it requires
      -- an extra wire to be added.
      clk_16MHz : in std_logic;

      -- All the control pins from the CPU socket
      cpu_PHI0_IN : in std_logic;
      cpu_PHI1_OUT : in std_logic;
      cpu_PHI2_OUT : in std_logic; -- best clock
      cpu_RDY : in std_logic;
      cpu_RnW : inout std_logic;
      cpu_SYNC : in std_logic;
      cpu_nIRQ : in std_logic;
      cpu_nNMI : in std_logic;
      cpu_nRESET : inout std_logic;
      cpu_nSO : in std_logic;

      -- General purpose pins, for passing clocks etc to the external device.
      -- ext_GP1, ext_GP3, and ext_GP4 are pulled up to 3V3, so should be used
      -- as active low chip enables for anything (driving the A/D bus, etc) that
      -- could have undesirable results during FPGA reprogramming or if the
      -- external device gets disconnected.
      ext_GP : inout std_logic_vector(12 downto 0) := (others => 'Z')

      -- GP0 convention: (is surrounded by ground plane) CPU clock; connected to
      -- cpu_PHI2_OUT.

      -- GP1 convention: (is surrounded by ground plane, has pullup to 3V3)
      -- global chip enable: 1=disable all buffers and shadowing, 0=enable
      -- buffer controls.  This is used to stop anything bad from happening
      -- while the external device is disconnected or tristated.

      -- GP2 convention: (is surrounded by ground plane) 16MHz clock; connected
      -- to clk_16MHz.

      -- GP3 convention: (has pullup to 3V3) /OE for data buffer.  When 1, the
      -- data buffer is disabled.  When 0, it's enabled.

      -- GP4 convention: (has pullup to 3V3) data buffer direction: 1=from CPU
      -- to connector, 0=from connector to CPU.

      -- GP5 convention: 1=onboard CPU, 0=external CPU. When 1, the address
      -- bus, RnW, SYNC, PHI1, and PHI2 are buffered from the CPU socket.
      -- When 0, all of these are buffered from the external connector (or
      -- PHI1/PHI2 are generated by the CPLD; not sure yet).

      -- GP6 convention: RnW
      -- GP7 convention: nRESET
      -- GP8 convention: RDY
      -- GP9 convention: /NMI
      -- GP10 convention: /IRQ
      -- GP11 convention:
      -- GP12 convention:

    );
end cpu_socket_expansion;

architecture Behavioural of cpu_socket_expansion is

  -- When '0', this disables all outputs and buffers

  signal global_enable : std_logic := '0';

  -- When '1', this forces A15:A13 = "110" (&C000-&DFFF address range), which
  -- will make the ULA think we're accessing the OS ROM.  If the (socketed)
  -- ROM is removed, this results in this tristating the data bus, letting the
  -- CPU access something without the ULA interfering.

  signal accessing_shadow_ram : std_logic := '0';

  -- When '1', this means the CPU is on the external connector (i.e. probably
  -- a soft-CPU implemented in an FPGA).  When '0', there is a 6502 plugged in
  -- to the onboard socket.

  signal cpu_is_external : std_logic := '0';

begin

  ext_GP(0) <= cpu_PHI2_OUT;

  global_enable <= not ext_GP(1);

  ext_GP(2) <= clk_16MHz;

  dbuf_nCE <= ext_GP(3) when global_enable = '1' else 'Z';
  dbuf_ext_to_cpu <= not ext_GP(4);

  cpu_is_external <= '0'; --not ext_GP(5);

  ext_GP(6) <= cpu_RnW when cpu_is_external = '0' else 'Z';
  cpu_RnW <= ext_GP(6) when cpu_is_external = '1' else 'Z';

  ext_GP(7) <= cpu_nRESET when cpu_is_external = '0' else 'Z';
  cpu_nRESET <= ext_GP(7) when cpu_is_external = '1' else 'Z';

  -- ABUF is always enabled
  abuf_nCE <= not global_enable;
  abuf_ext_to_cpu <= cpu_is_external;

  -- Buffer A15:13 from socketed CPU (or external CPU via ABUFH) to motherboard
  cpu_A15_1 <= '1' when accessing_shadow_ram = '1' else cpu_A15_2;
  cpu_A14_1 <= '1' when accessing_shadow_ram = '1' else cpu_A14_2;
  cpu_A13_1 <= '0' when accessing_shadow_ram = '1' else cpu_A13_2;

end Behavioural;
